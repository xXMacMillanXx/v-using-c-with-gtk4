module graphene

#flag -I/usr/include/graphene-1.0 -L/usr/lib64
#flag -I/lib64/graphene-1.0/include -L/usr/lib64
#flag -lgraphene-1.0