module pango

#flag -I/usr/include/pango-1.0 -L/usr/lib64
#flag -lpango-1.0