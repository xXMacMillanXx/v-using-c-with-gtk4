module harfbuzz

#flag -I/usr/include/harfbuzz -L/usr/lib64
#flag -lharfbuzz